-- Confics specific for fast poly_fir

package bench_config is
    constant USE_SLOW_POLY_FIR : boolean := false;

    constant STROBE_DATA_DELAY : natural := 2;
end;
