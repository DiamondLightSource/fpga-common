-- Confics specific for slow poly_fir

package bench_config is
    constant USE_SLOW_POLY_FIR : boolean := true;

    constant STROBE_DATA_DELAY : natural := 20;
end;
