../../common/sim_support.vhd